version https://git-lfs.github.com/spec/v1
oid sha256:9520618d55c475062ef8cb19008b39b24fc4c2544681b9a6012c09d13afc3195
size 663
